// Inverter
module inverter(
input a,
output x);

assign x = ~a;
endmodule
